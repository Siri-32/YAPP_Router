/*-------------------------------------------------------------------------
File name   : router.svh
Title       : Module UVC Files
----------------------------------------------------------------------*/

`include "router_scoreboard.sv"
`include "router_reference.sv"
`include "router_module_env.sv"
